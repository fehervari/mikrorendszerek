//******************************************************************************
//* Verilog functions used in the memory controller.                           *
//*                                                                            *
//* Written by   : Tamas Raikovich                                             *
//* Version      : 2.0                                                         *
//* Last modified: 2012.10.21.                                                 *
//******************************************************************************


//******************************************************************************
//* Base 2 logarithm function.                                                 *
//******************************************************************************
function integer log2(input integer x);
   for (log2 = 0; x > 0; log2 = log2 + 1)
      x = x >> 1;
endfunction
